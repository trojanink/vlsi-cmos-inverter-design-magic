magic
tech scmos
timestamp 1477900137
<< nwell >>
rect -42 52 -6 74
<< polysilicon >>
rect -37 61 -35 63
rect -29 61 -27 63
rect -21 61 -19 63
rect -13 61 -11 63
rect -37 40 -35 58
rect -29 40 -27 58
rect -21 40 -19 58
rect -13 40 -11 58
rect -37 35 -35 37
rect -29 35 -27 37
rect -21 35 -19 37
rect -13 35 -11 37
<< ndiffusion >>
rect -38 37 -37 40
rect -35 37 -34 40
rect -30 37 -29 40
rect -27 37 -26 40
rect -22 37 -21 40
rect -19 37 -18 40
rect -14 37 -13 40
rect -11 37 -10 40
<< pdiffusion >>
rect -38 58 -37 61
rect -35 58 -34 61
rect -30 58 -29 61
rect -27 58 -26 61
rect -22 58 -21 61
rect -19 58 -18 61
rect -14 58 -13 61
rect -11 58 -10 61
<< metal1 >>
rect -38 72 -34 76
rect -30 72 -26 76
rect -22 72 -18 76
rect -14 72 -10 76
rect -34 62 -30 72
rect -42 53 -38 58
rect -10 53 -6 58
rect -46 50 -2 53
rect -42 41 -38 50
rect -34 44 -14 47
rect -34 41 -30 44
rect -18 41 -14 44
rect -26 33 -22 37
rect -10 33 -6 37
rect -38 29 -34 33
rect -30 29 -26 33
rect -22 29 -18 33
rect -14 29 -10 33
<< ntransistor >>
rect -37 37 -35 40
rect -29 37 -27 40
rect -21 37 -19 40
rect -13 37 -11 40
<< ptransistor >>
rect -37 58 -35 61
rect -29 58 -27 61
rect -21 58 -19 61
rect -13 58 -11 61
<< ndcontact >>
rect -42 37 -38 41
rect -34 37 -30 41
rect -26 37 -22 41
rect -18 37 -14 41
rect -10 37 -6 41
<< pdcontact >>
rect -42 58 -38 62
rect -34 58 -30 62
rect -26 58 -22 62
rect -18 58 -14 62
rect -10 58 -6 62
<< nbccdiffcontact >>
rect -34 72 -30 76
<< psubstratepcontact >>
rect -42 29 -38 33
rect -34 29 -30 33
rect -26 29 -22 33
rect -18 29 -14 33
rect -10 29 -6 33
<< nsubstratencontact >>
rect -42 72 -38 76
rect -26 72 -22 76
rect -18 72 -14 76
rect -10 72 -6 76
<< labels >>
rlabel metal1 -6 51 -2 51 7 out
rlabel metal1 -46 51 -42 51 3 in
rlabel metal1 -30 74 -26 74 5 vdd
rlabel metal1 -29 31 -25 31 1 gnd
rlabel polysilicon -37 61 -35 63 1 b
rlabel polysilicon -29 61 -27 63 1 a
rlabel polysilicon -21 61 -19 63 1 c
rlabel polysilicon -13 61 -11 63 1 d
<< end >>
